module initial_permutation (output_text, plain_text);

input [64:1] plain_text;
output wire [64:1] output_text;

assign output_text[1] = plain_text[58];
assign output_text[2] = plain_text[50];
assign output_text[3] = plain_text[42];
assign output_text[4] = plain_text[34];
assign output_text[5] = plain_text[26];
assign output_text[6] = plain_text[18];
assign output_text[7] = plain_text[10];
assign output_text[8] = plain_text[2];
assign output_text[9] = plain_text[60];
assign output_text[10] = plain_text[52];
assign output_text[11] = plain_text[44];
assign output_text[12] = plain_text[36];
assign output_text[13] = plain_text[28];
assign output_text[14] = plain_text[20];
assign output_text[15] = plain_text[12];
assign output_text[16] = plain_text[4];
assign output_text[17] = plain_text[62];
assign output_text[18] = plain_text[54];
assign output_text[19] = plain_text[46];
assign output_text[20] = plain_text[38];
assign output_text[21] = plain_text[30];
assign output_text[22] = plain_text[22];
assign output_text[23] = plain_text[14];
assign output_text[24] = plain_text[6];
assign output_text[25] = plain_text[64];
assign output_text[26] = plain_text[56];
assign output_text[27] = plain_text[48];
assign output_text[28] = plain_text[40];
assign output_text[29] = plain_text[32];
assign output_text[30] = plain_text[24];
assign output_text[31] = plain_text[16];
assign output_text[32] = plain_text[8];
assign output_text[33] = plain_text[57];
assign output_text[34] = plain_text[49];
assign output_text[35] = plain_text[41];
assign output_text[36] = plain_text[33];
assign output_text[37] = plain_text[25];
assign output_text[38] = plain_text[17];
assign output_text[39] = plain_text[9];
assign output_text[40] = plain_text[1];
assign output_text[41] = plain_text[59];
assign output_text[42] = plain_text[51];
assign output_text[43] = plain_text[43];
assign output_text[44] = plain_text[35];
assign output_text[45] = plain_text[27];
assign output_text[46] = plain_text[19];
assign output_text[47] = plain_text[11];
assign output_text[48] = plain_text[3];
assign output_text[49] = plain_text[61];
assign output_text[50] = plain_text[53];
assign output_text[51] = plain_text[45];
assign output_text[52] = plain_text[37];
assign output_text[53] = plain_text[29];
assign output_text[54] = plain_text[21];
assign output_text[55] = plain_text[13];
assign output_text[56] = plain_text[5];
assign output_text[57] = plain_text[63];
assign output_text[58] = plain_text[55];
assign output_text[59] = plain_text[47];
assign output_text[60] = plain_text[39];
assign output_text[61] = plain_text[31];
assign output_text[62] = plain_text[23];
assign output_text[63] = plain_text[15];
assign output_text[64] = plain_text[7];

endmodule