module final_permutation (cipher_text, input_text);

input [64:1] input_text;
output reg [64:1] cipher_text;

assign cipher_text[1] = input_text[40];
assign cipher_text[2] = input_text[8];
assign cipher_text[3] = input_text[48];
assign cipher_text[4] = input_text[16];
assign cipher_text[5] = input_text[56];
assign cipher_text[6] = input_text[24];
assign cipher_text[7] = input_text[64];
assign cipher_text[8] = input_text[32];
assign cipher_text[9] = input_text[39];
assign cipher_text[10] = input_text[7];
assign cipher_text[11] = input_text[47];
assign cipher_text[12] = input_text[15];
assign cipher_text[13] = input_text[55];
assign cipher_text[14] = input_text[23];
assign cipher_text[15] = input_text[63];
assign cipher_text[16] = input_text[31];
assign cipher_text[17] = input_text[38];
assign cipher_text[18] = input_text[6];
assign cipher_text[19] = input_text[46];
assign cipher_text[20] = input_text[14];
assign cipher_text[21] = input_text[54];
assign cipher_text[22] = input_text[22];
assign cipher_text[23] = input_text[62];
assign cipher_text[24] = input_text[30];
assign cipher_text[25] = input_text[37];
assign cipher_text[26] = input_text[5];
assign cipher_text[27] = input_text[45];
assign cipher_text[28] = input_text[13];
assign cipher_text[29] = input_text[53];
assign cipher_text[30] = input_text[21];
assign cipher_text[31] = input_text[61];
assign cipher_text[32] = input_text[29];
assign cipher_text[33] = input_text[36];
assign cipher_text[34] = input_text[4];
assign cipher_text[35] = input_text[44];
assign cipher_text[36] = input_text[12];
assign cipher_text[37] = input_text[52];
assign cipher_text[38] = input_text[20];
assign cipher_text[39] = input_text[60];
assign cipher_text[40] = input_text[28];
assign cipher_text[41] = input_text[35];
assign cipher_text[42] = input_text[3];
assign cipher_text[43] = input_text[43];
assign cipher_text[44] = input_text[11];
assign cipher_text[45] = input_text[51];
assign cipher_text[46] = input_text[19];
assign cipher_text[47] = input_text[59];
assign cipher_text[48] = input_text[27];
assign cipher_text[49] = input_text[34];
assign cipher_text[50] = input_text[2];
assign cipher_text[51] = input_text[42];
assign cipher_text[52] = input_text[10];
assign cipher_text[53] = input_text[50];
assign cipher_text[54] = input_text[18];
assign cipher_text[55] = input_text[58];
assign cipher_text[56] = input_text[26];
assign cipher_text[57] = input_text[33];
assign cipher_text[58] = input_text[1];
assign cipher_text[59] = input_text[41];
assign cipher_text[60] = input_text[9];
assign cipher_text[61] = input_text[49];
assign cipher_text[62] = input_text[17];
assign cipher_text[63] = input_text[57];
assign cipher_text[64] = input_text[25];

endmodule