module permutation_choice_one (perm_choice_one_output, perm_choice_one_input);

input [64:1] perm_choice_one_input;
output [56:1] perm_choice_one_output;

assign perm_choice_one_output[1] = perm_choice_one_input[57];
assign perm_choice_one_output[2] = perm_choice_one_input[49];
assign perm_choice_one_output[3] = perm_choice_one_input[41];
assign perm_choice_one_output[4] = perm_choice_one_input[33];
assign perm_choice_one_output[5] = perm_choice_one_input[25];
assign perm_choice_one_output[6] = perm_choice_one_input[17];
assign perm_choice_one_output[7] = perm_choice_one_input[9];
assign perm_choice_one_output[8] = perm_choice_one_input[1];
assign perm_choice_one_output[9] = perm_choice_one_input[58];
assign perm_choice_one_output[10] = perm_choice_one_input[50];
assign perm_choice_one_output[11] = perm_choice_one_input[42];
assign perm_choice_one_output[12] = perm_choice_one_input[34];
assign perm_choice_one_output[13] = perm_choice_one_input[26];
assign perm_choice_one_output[14] = perm_choice_one_input[18];
assign perm_choice_one_output[15] = perm_choice_one_input[10];
assign perm_choice_one_output[16] = perm_choice_one_input[2];
assign perm_choice_one_output[17] = perm_choice_one_input[59];
assign perm_choice_one_output[18] = perm_choice_one_input[51];
assign perm_choice_one_output[19] = perm_choice_one_input[43];
assign perm_choice_one_output[20] = perm_choice_one_input[35];
assign perm_choice_one_output[21] = perm_choice_one_input[27];
assign perm_choice_one_output[22] = perm_choice_one_input[19];
assign perm_choice_one_output[23] = perm_choice_one_input[11];
assign perm_choice_one_output[24] = perm_choice_one_input[3];
assign perm_choice_one_output[25] = perm_choice_one_input[60];
assign perm_choice_one_output[26] = perm_choice_one_input[52];
assign perm_choice_one_output[27] = perm_choice_one_input[44];
assign perm_choice_one_output[28] = perm_choice_one_input[36];
assign perm_choice_one_output[29] = perm_choice_one_input[63];
assign perm_choice_one_output[30] = perm_choice_one_input[55];
assign perm_choice_one_output[31] = perm_choice_one_input[47];
assign perm_choice_one_output[32] = perm_choice_one_input[39];
assign perm_choice_one_output[33] = perm_choice_one_input[31];
assign perm_choice_one_output[34] = perm_choice_one_input[23];
assign perm_choice_one_output[35] = perm_choice_one_input[15];
assign perm_choice_one_output[36] = perm_choice_one_input[7];
assign perm_choice_one_output[37] = perm_choice_one_input[62];
assign perm_choice_one_output[38] = perm_choice_one_input[55];
assign perm_choice_one_output[39] = perm_choice_one_input[46];
assign perm_choice_one_output[40] = perm_choice_one_input[38];
assign perm_choice_one_output[41] = perm_choice_one_input[30];
assign perm_choice_one_output[42] = perm_choice_one_input[22];
assign perm_choice_one_output[43] = perm_choice_one_input[14];
assign perm_choice_one_output[44] = perm_choice_one_input[6];
assign perm_choice_one_output[45] = perm_choice_one_input[61];
assign perm_choice_one_output[46] = perm_choice_one_input[53];
assign perm_choice_one_output[47] = perm_choice_one_input[45];
assign perm_choice_one_output[48] = perm_choice_one_input[37];
assign perm_choice_one_output[49] = perm_choice_one_input[29];
assign perm_choice_one_output[50] = perm_choice_one_input[21];
assign perm_choice_one_output[51] = perm_choice_one_input[13];
assign perm_choice_one_output[52] = perm_choice_one_input[5];
assign perm_choice_one_output[53] = perm_choice_one_input[28];
assign perm_choice_one_output[54] = perm_choice_one_input[20];
assign perm_choice_one_output[55] = perm_choice_one_input[12];
assign perm_choice_one_output[56] = perm_choice_one_input[4];

endmodule